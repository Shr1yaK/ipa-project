module pc(
    input clk,
)
endmodule